`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UT ECE
// Engineer: Jan C. Rubio
// UT EID: jcr4698
// 
// Create Date: 11/21/2021 11:12:38 PM
// Design Name: Stopwatch/Timer
// Module Name: stopwatch_state_machine
// Project Name: Lab 6
// Target Devices: Basys3
// Description: State machine of programmable stopwatch/timer with RTL Design.
// 
//////////////////////////////////////////////////////////////////////////////////


module stopwatch_state_machine(
    input clk,
    input [6:0] in0,
    input [6:0] in1,
    input [6:0] in2,
    input [6:0] in3,
    output reg [3:0] an,
    output reg [6:0] sseg
    );
    
    // TODO: state machine logic for 7 segment display
    
    // TODO: state machine logic for data path
    
endmodule
