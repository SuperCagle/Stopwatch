`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UT ECE
// Engineer: Jan C. Rubio
// UT EID: jcr4698
// 
// Create Date: 11/21/2021 11:12:38 PM
// Design Name: Stopwatch/Timer
// Module Name: upCount
// Project Name: Lab 6
// Target Devices: Basys3
// Description:  Up counter with optional initial time programmable stopwatch/timer. 
// Design will be implemented using RTL-design methodology with 4 modes.
// 
//////////////////////////////////////////////////////////////////////////////////


module upCount(
    input clk,
    input setTime,
    input stop,
    input clr,
    input di0,
    input di1,
    input di2,
    input di3
    );
    
    // TODO: timer down implementation
    
endmodule
