`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UT ECE
// Engineer: Jan C. Rubio
// UT EID: jcr4698
// 
// Create Date: 11/21/2021 11:12:38 PM
// Design Name: Stopwatch/Timer
// Module Name: stopwatch_state_machine
// Project Name: Lab 6
// Target Devices: Basys3
// Description:  programmable stopwatch/timer design will be implemented using 
// RTL-design methodology with 4 modes.
// 
//////////////////////////////////////////////////////////////////////////////////


module time_mux_state_machine(

    );
endmodule
